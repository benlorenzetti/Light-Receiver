*** stage2.cir ***

Vcc cc gnd DC 5

************************** Stage I Equivalent *******************
Vmirror mirror gnd DC 1
Vin out1 gnd 1m AC 1 PULSE (0 1m 0 1n 1n 50n 100n)
Rc1 out1 in2 100

************************* Stage II ******************************
R5 cc b7 2.74k
Re5 e5 gnd 342
Re6 e6 gnd 25
R7 cc b8 666
R8 b8 gnd 2000
Ce7 e7 gnd 100u IC=1
C5 n5 b7 100n
L5 in2 n5 1u

Q5 b7 mirror e5 n3904
Q6 e7 mirror e6 n3904
Q7 c7 b7 e7 n2369
Q8 cc b8 b9 n3904
Q9 c9 b9 c7 n2369

*** Capacitative Coupling to Stage III ***
Rdif cc c9 100
Cload c9 out2p 10u
Rload out2p gnd 100k
*** Transformer Coupling to Stage III ****
*X1 cc c9 out2p gnd murata76615
*Rdif out2p gnd 100

.subckt murata76615 1 2 3 4
Lleakp 1 11 2u
Rp 11 111 1.00
Lp 111 2 3200u
Lleaks 3 33 2u
Rs 33 333 1.00
Ls 333 4 3200u
K Lp Ls 1
.ends murata76615

.model n3904 npn (IS=1E-14 VAF=100 Bf=300 IKF=0.4 XTB=1.5 BR=4 CJC=4E-12 CJE=8E-12 RB=20 RC=0.1 RE=0.1 TR=250E-9 TF=350E-12 ITF=1 VTF=2 XTF=3 Vceo=40 Icrating=200m)
.model n2369 npn (Is=44.14f Xti=3 Eg=1.11 Vaf=100 Bf=78.32 Ne=1.389 Ise=91.95f Ikf=.3498 Xtb=1.5 Br=12.69m Nc=2 Isc=0 Ikr=0 Rc=.6 Cjc=2.83p Mjc=86.19m Vjc=.75 Fc=.5 Cje=4.5p Mje=.2418 Vje=.75 Tr=1.073u Tf=227.6p Itf=.3 Vtf=4 Xtf=4 Rb=10 Vceo=15 Icrating=200m)

.control
ac dec 100 1 100G
plot vdb(out2p)
plot vp(out2p)
wrdata spice2 vdb(out2p) vp(out2p)
tran 0.1ns 1000ns
plot v(out1)
plot v(out2p)

