*** transimpedance.cir ***

Vcc cc gnd DC 5

Isigma in gnd AC 1 SIN (0 1 10Meg)
Csigma in gnd 960p

Re0 me0 gnd 100
Re1 me1 gnd 10
R0 cc mirror 2.4k
R1 cc b1 414
R2 b1 gnd 276
Rc cc out 90
Rl out gnd 100k

Q1 out b1 in model2n3904
Qm1 in mirror me1 model2n3904
Qm0 mirror mirror me0 model2n3904

.model model2n3904 npn (bf=100 vaf=200 cje=18p cjc=4p)

.control
op
ac dec 100 100k 1000Meg
plot vdb(out)
plot vp(out)
wrdata spice-output vdb(out) vp(out)
.end
