*** ./s2-BJT-d3 ***
*f3=10000000000, f4=100, f5=1000, f6=100000
Vcc cc gnd DC 5
Vc1 indc gnd DC 3.075000
Vin in indc 1m AC 1 SIN (0 1 10Meg)
Vmirror mirror gnd DC 1.016000
Rc1 c1 in 250.000000
L6 c1 n5 147.269162n
R5 n5 b3 17.109156k
C5 n5 b3 17200.000000n
R7 cc b4 63.156723
R8 b4 gnd 107.537124
Rc4 cc out 250.669035
Re3 me3 gnd 26.419721
Ce3 e3 gnd 9.302326u

Q3 c3 b3 e3 2n3904
Qm3 e3 mirror me3 2n3904
Q4 out b4 c3 2n3904
.model 2n3904 npn (bf=100.000000 vaf=200 cje=18p cjc=4p)
.control
ac dec 100 10 1000Meg
plot vdb(out)
plot vp(out)
wrdata spice-output vdb(out) vp(out)
