*** CE-Amplifier.cir ***
*
Vcc cc gnd DC 5
Vinput in inac 1m AC 1 SIN (0 1 10Meg)

.param q3beta=100.000000
Vc1 in gnd DC 3.075000
Vmirror mirror gnd DC 1.016000
Rc1 inac c1 250.000000
R4 c1 b3 107.250000k
C4 c1 b3 148051.109853p
Rc3 cc out 1575.000000
Re3 me3 gnd 166.000000
Ce3 e3 gnd 1.480511u
R5 b4 cc 396.825397
R6 b4 gnd 675.675676


Q3 c3 b3 e3 model2n3904
Qm3 e3 mirror me3 model2n3904
Q4 out b4 c3 model2n3904

.model model2n3904 npn (bf={q3beta} vaf=200 cje=18p cjc=0.4p)

.control
ac dec 100 100 1000Meg
plot vdb(out)
plot vp(out)
wrdata spice-output vdb(out) vp(out)
