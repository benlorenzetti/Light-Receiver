*** transimpedance.cir ***

Vcc cc gnd DC 5

Isigma in gnd DC 1u AC 1 SIN (0 200n 10Meg)
Csigma in gnd 960p

Re1 me1 gnd 10
Re2 me2 cc 10
Rc out cc 250
R0 b2 mirror 1906
R1 e0 gnd 100
R2 b2 cc 745
R3 cc b1 92.5
R4 b1 gnd 69.8

Q0 mirror mirror e0 model2n3904
Q1 out b1 in model2n3904
Qm1 in mirror me1 model2n3904
Q2 out b2 e2 model2n3906

.model model2n3904 npn (bf=100 vaf=200 cje=18p cjc=4p)
.model model2n3906 pnp (bf=100 vaf=200 cje=25p cjc=6p)

.control
op
ac dec 100 100k 1000Meg
plot vdb(out)
plot vp(out)
wrdata spice-output vdb(out) vp(out)
.end
