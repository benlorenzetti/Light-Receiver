*** stage1.cir ***

Vcc cc gnd DC 5

Iamb in gnd DC 1u
Iin in gnd 1m AC 1 SIN (0 1 10Meg)
Csigma in gnd 15p

R0 cc mirror 1.7k
R1 cc b2 723
R2 b2 gnd 884
R3 e3 gnd 10.6
R4 e4 gnd 106

Rc1 cc out1 100

Q1 out1 b1 in n2369
Q2 cc b2 b1 n3904
Q3 in mirror e3 n3904
Q4 mirror mirror e4 n3904

.model n3904 npn (IS=1E-14 VAF=100 Bf=300 IKF=0.4 XTB=1.5 BR=4 CJC=4E-12 CJE=8E-12 RB=20 RC=0.1 RE=0.1 TR=250E-9 TF=350E-12 ITF=1 VTF=2 XTF=3 Vceo=40 Icrating=200m)
.model n2369 npn (Is=44.14f Xti=3 Eg=1.11 Vaf=100 Bf=78.32 Ne=1.389 Ise=91.95f Ikf=.3498 Xtb=1.5 Br=12.69m Nc=2 Isc=0 Ikr=0 Rc=.6 Cjc=2.83p Mjc=86.19m Vjc=.75 Fc=.5 Cje=4.5p Mje=.2418 Vje=.75 Tr=1.073u Tf=227.6p Itf=.3 Vtf=4 Xtf=4 Rb=10 Vceo=15 Icrating=200m)

.control
ac dec 100 1 100G
plot vdb(out1)
plot vp(out1)
wrdata spice1 vdb(out1) vp(out1)
